class stimulus;
	//rand reg [3:0] address;
	//rand reg [3:0] address2;
	//rand reg [3:0] address3;
	//rand reg [3:0] address4;
	//rand reg [3:0] address5;
	//rand reg [3:0] address6;
	//rand reg [3:0] address7;
	//rand reg [3:0] address8;

	rand reg [15:0] din;
	rand reg [2:0]count;
endclass
