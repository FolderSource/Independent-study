   class scoreboardt;
      reg [7:0] store;
      reg [7:0] var_x;
      reg [7:0] var_z;
      //reg [7:0] counter1;
      //reg [7:0] counter2;
      //reg [7:0] array1[10:0];
      //array1.push_front(0);
      //reg[7:0] array1[$];
      reg digit_clk;
      reg dout_flag;
      //reg [7:0] array2[9999:0];
   endclass
